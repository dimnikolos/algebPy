-- Top Level Structural Model for MIPS Processor Core
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY TEST IS
END TEST;
ARCHITECTURE BEH OF TEST IS
COMPONENT MIPS PORT (clock : IN STD_LOGIC;
	reset : IN STD_LOGIC);
END COMPONENT;

COMPONENT THECLOCK PORT (clock: OUT STD_LOGIC; reset: OUT STD_LOGIC);
END COMPONENT;

SIGNAL CLK: STD_LOGIC;
SIGNAL RST: STD_LOGIC;
BEGIN

PROC: MIPS PORT MAP(
	clock => CLK,
	reset => RST);
CLKGEN: THECLOCK PORT MAP(
	clock => CLK,
	reset => RST);
END BEH;

